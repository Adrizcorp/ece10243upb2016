module mux_nco_freq(
		input [2:0]sel,
		output [31:0]out
	);

assign out[31:0]=(sel[2:0]==3'd0)	?  32'd85:
				     (sel[2:0]==3'd1)	?	32'd12887:
					  (sel[2:0]==3'd2)	?	32'd171799:
					  (sel[2:0]==3'd3)	?	32'd429497:
					  (sel[2:0]==3'd4)	?	32'd687195:
					  (sel[2:0]==3'd5)	?	32'd773095:
					  (sel[2:0]==3'd6)	?	32'd858994:
					  32'd1717987;
/*	
85   //1 Hz 
12887  //150 Hz
171799 //2000 Hz
429497 //5000 Hz
687195 //8000 Hz
773095 //9000 Hz
858994 //10000 Hz
1717987//200000
*/
	
endmodule
