// nios_practica.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module nios_practica (
		input  wire        clk_clk,            //         clk.clk
		output wire [31:0] div_freq_export,    //    div_freq.export
		output wire [7:0]  leds_export,        //        leds.export
		output wire [15:0] noise_export,       //       noise.export
		output wire        noise_en_export,    //    noise_en.export
		output wire        noise_pulse_export, // noise_pulse.export
		input  wire        reset_reset_n,      //       reset.reset_n
		output wire [9:0]  sel_nota_export,    //    sel_nota.export
		input  wire [3:0]  sw_export,          //          sw.export
		output wire        timer_export,       //       timer.export
		input  wire        uart_rxd,           //        uart.rxd
		output wire        uart_txd            //            .txd
	);

	wire         pll_outclk0_clk;                                                     // pll:outclk_0 -> [RAM_jesus:clk, cpu:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, rst_controller:clk, rst_controller_002:clk, uart:clk]
	wire  [31:0] cpu_data_master_readdata;                                            // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                         // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                         // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                                             // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                          // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                               // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                           // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                     // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                  // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                                      // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                         // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;              // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;           // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_chipselect; // mm_interconnect_0:timer_ece10243upb2016_0_avalon_slave_0_chipselect -> timer_ece10243upb2016_0:timer_chipselect
	wire  [31:0] mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_readdata;   // timer_ece10243upb2016_0:timer_readdata -> mm_interconnect_0:timer_ece10243upb2016_0_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_address;    // mm_interconnect_0:timer_ece10243upb2016_0_avalon_slave_0_address -> timer_ece10243upb2016_0:timer_address
	wire         mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_write;      // mm_interconnect_0:timer_ece10243upb2016_0_avalon_slave_0_write -> timer_ece10243upb2016_0:timer_write
	wire  [31:0] mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_writedata;  // mm_interconnect_0:timer_ece10243upb2016_0_avalon_slave_0_writedata -> timer_ece10243upb2016_0:timer_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                      // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                   // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                   // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                       // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                          // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                    // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                         // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                     // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_jesus_s1_chipselect;                           // mm_interconnect_0:RAM_jesus_s1_chipselect -> RAM_jesus:chipselect
	wire  [31:0] mm_interconnect_0_ram_jesus_s1_readdata;                             // RAM_jesus:readdata -> mm_interconnect_0:RAM_jesus_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_jesus_s1_address;                              // mm_interconnect_0:RAM_jesus_s1_address -> RAM_jesus:address
	wire   [3:0] mm_interconnect_0_ram_jesus_s1_byteenable;                           // mm_interconnect_0:RAM_jesus_s1_byteenable -> RAM_jesus:byteenable
	wire         mm_interconnect_0_ram_jesus_s1_write;                                // mm_interconnect_0:RAM_jesus_s1_write -> RAM_jesus:write
	wire  [31:0] mm_interconnect_0_ram_jesus_s1_writedata;                            // mm_interconnect_0:RAM_jesus_s1_writedata -> RAM_jesus:writedata
	wire         mm_interconnect_0_ram_jesus_s1_clken;                                // mm_interconnect_0:RAM_jesus_s1_clken -> RAM_jesus:clken
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                    // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                                     // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                  // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                   // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                     // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                 // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                                // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                                  // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                                   // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                                      // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                             // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                                     // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                                 // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_div_freq_s1_chipselect;                            // mm_interconnect_0:div_freq_s1_chipselect -> div_freq:chipselect
	wire  [31:0] mm_interconnect_0_div_freq_s1_readdata;                              // div_freq:readdata -> mm_interconnect_0:div_freq_s1_readdata
	wire   [1:0] mm_interconnect_0_div_freq_s1_address;                               // mm_interconnect_0:div_freq_s1_address -> div_freq:address
	wire         mm_interconnect_0_div_freq_s1_write;                                 // mm_interconnect_0:div_freq_s1_write -> div_freq:write_n
	wire  [31:0] mm_interconnect_0_div_freq_s1_writedata;                             // mm_interconnect_0:div_freq_s1_writedata -> div_freq:writedata
	wire         mm_interconnect_0_sys_clk_s1_chipselect;                             // mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_s1_readdata;                               // sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_s1_address;                                // mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	wire         mm_interconnect_0_sys_clk_s1_write;                                  // mm_interconnect_0:sys_clk_s1_write -> sys_clk:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_s1_writedata;                              // mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	wire         mm_interconnect_0_noise_s1_chipselect;                               // mm_interconnect_0:noise_s1_chipselect -> noise:chipselect
	wire  [31:0] mm_interconnect_0_noise_s1_readdata;                                 // noise:readdata -> mm_interconnect_0:noise_s1_readdata
	wire   [1:0] mm_interconnect_0_noise_s1_address;                                  // mm_interconnect_0:noise_s1_address -> noise:address
	wire         mm_interconnect_0_noise_s1_write;                                    // mm_interconnect_0:noise_s1_write -> noise:write_n
	wire  [31:0] mm_interconnect_0_noise_s1_writedata;                                // mm_interconnect_0:noise_s1_writedata -> noise:writedata
	wire         mm_interconnect_0_noise_en_s1_chipselect;                            // mm_interconnect_0:noise_en_s1_chipselect -> noise_en:chipselect
	wire  [31:0] mm_interconnect_0_noise_en_s1_readdata;                              // noise_en:readdata -> mm_interconnect_0:noise_en_s1_readdata
	wire   [1:0] mm_interconnect_0_noise_en_s1_address;                               // mm_interconnect_0:noise_en_s1_address -> noise_en:address
	wire         mm_interconnect_0_noise_en_s1_write;                                 // mm_interconnect_0:noise_en_s1_write -> noise_en:write_n
	wire  [31:0] mm_interconnect_0_noise_en_s1_writedata;                             // mm_interconnect_0:noise_en_s1_writedata -> noise_en:writedata
	wire         mm_interconnect_0_sel_nota_s1_chipselect;                            // mm_interconnect_0:sel_nota_s1_chipselect -> sel_nota:chipselect
	wire  [31:0] mm_interconnect_0_sel_nota_s1_readdata;                              // sel_nota:readdata -> mm_interconnect_0:sel_nota_s1_readdata
	wire   [1:0] mm_interconnect_0_sel_nota_s1_address;                               // mm_interconnect_0:sel_nota_s1_address -> sel_nota:address
	wire         mm_interconnect_0_sel_nota_s1_write;                                 // mm_interconnect_0:sel_nota_s1_write -> sel_nota:write_n
	wire  [31:0] mm_interconnect_0_sel_nota_s1_writedata;                             // mm_interconnect_0:sel_nota_s1_writedata -> sel_nota:writedata
	wire         mm_interconnect_0_noise_pulse_s1_chipselect;                         // mm_interconnect_0:noise_pulse_s1_chipselect -> noise_pulse:chipselect
	wire  [31:0] mm_interconnect_0_noise_pulse_s1_readdata;                           // noise_pulse:readdata -> mm_interconnect_0:noise_pulse_s1_readdata
	wire   [1:0] mm_interconnect_0_noise_pulse_s1_address;                            // mm_interconnect_0:noise_pulse_s1_address -> noise_pulse:address
	wire         mm_interconnect_0_noise_pulse_s1_write;                              // mm_interconnect_0:noise_pulse_s1_write -> noise_pulse:write_n
	wire  [31:0] mm_interconnect_0_noise_pulse_s1_writedata;                          // mm_interconnect_0:noise_pulse_s1_writedata -> noise_pulse:writedata
	wire         irq_mapper_receiver1_irq;                                            // uart:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                                            // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                                         // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver0_irq;                                            // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                       // timer_ece10243upb2016_0:timer_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                            // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                   // sys_clk:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [RAM_jesus:reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [RAM_jesus:reset_req, cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                       // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [div_freq:reset_n, irq_synchronizer_001:receiver_reset, leds:reset_n, mm_interconnect_0:sw_reset_reset_bridge_in_reset_reset, sw:reset_n, sys_clk:reset_n]
	wire         rst_controller_002_reset_out_reset;                                  // rst_controller_002:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                  // rst_controller_003:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:timer_ece10243upb2016_0_reset_reset_bridge_in_reset_reset, noise:reset_n, noise_en:reset_n, noise_pulse:reset_n, sel_nota:reset_n, timer_ece10243upb2016_0:reset]

	nios_practica_RAM_jesus ram_jesus (
		.clk        (pll_outclk0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_ram_jesus_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_jesus_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_jesus_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_jesus_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_jesus_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_jesus_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_jesus_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)         //       .reset_req
	);

	nios_practica_cpu cpu (
		.clk                                 (pll_outclk0_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios_practica_div_freq div_freq (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_div_freq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_div_freq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_div_freq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_div_freq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_div_freq_s1_readdata),   //                    .readdata
		.out_port   (div_freq_export)                           // external_connection.export
	);

	nios_practica_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	nios_practica_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	nios_practica_noise noise (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_noise_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_noise_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_noise_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_noise_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_noise_s1_readdata),   //                    .readdata
		.out_port   (noise_export)                           // external_connection.export
	);

	nios_practica_noise_en noise_en (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_noise_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_noise_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_noise_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_noise_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_noise_en_s1_readdata),   //                    .readdata
		.out_port   (noise_en_export)                           // external_connection.export
	);

	nios_practica_noise_en noise_pulse (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_noise_pulse_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_noise_pulse_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_noise_pulse_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_noise_pulse_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_noise_pulse_s1_readdata),   //                    .readdata
		.out_port   (noise_pulse_export)                           // external_connection.export
	);

	nios_practica_pll pll (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.locked   ()                 //  locked.export
	);

	nios_practica_sel_nota sel_nota (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_sel_nota_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sel_nota_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sel_nota_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sel_nota_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sel_nota_s1_readdata),   //                    .readdata
		.out_port   (sel_nota_export)                           // external_connection.export
	);

	nios_practica_sw sw (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata),    //                    .readdata
		.in_port  (sw_export)                            // external_connection.export
	);

	nios_practica_sys_clk sys_clk (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)        //   irq.irq
	);

	nios_practica_timer_ece10243upb2016_0 timer_ece10243upb2016_0 (
		.clk              (clk_clk),                                                             //          clock.clk
		.timer_address    (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_address),    // avalon_slave_0.address
		.timer_chipselect (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_chipselect), //               .chipselect
		.timer_readdata   (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_readdata),   //               .readdata
		.timer_write      (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_write),      //               .write
		.timer_writedata  (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_writedata),  //               .writedata
		.reset            (rst_controller_003_reset_out_reset),                                  //          reset.reset
		.toggle           (timer_export),                                                        //          timer.export
		.timer_irq        (irq_synchronizer_receiver_irq)                                        //      interrupt.irq
	);

	nios_practica_uart uart (
		.clk           (pll_outclk0_clk),                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	nios_practica_mm_interconnect_0 mm_interconnect_0 (
		.clk_50mhz_clk_clk                                         (clk_clk),                                                             //                                       clk_50mhz_clk.clk
		.pll_outclk0_clk                                           (pll_outclk0_clk),                                                     //                                         pll_outclk0.clk
		.cpu_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                                      //                     cpu_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset               (rst_controller_002_reset_out_reset),                                  //               jtag_uart_reset_reset_bridge_in_reset.reset
		.sw_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),                                  //                      sw_reset_reset_bridge_in_reset.reset
		.timer_ece10243upb2016_0_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                                  // timer_ece10243upb2016_0_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                   (cpu_data_master_address),                                             //                                     cpu_data_master.address
		.cpu_data_master_waitrequest                               (cpu_data_master_waitrequest),                                         //                                                    .waitrequest
		.cpu_data_master_byteenable                                (cpu_data_master_byteenable),                                          //                                                    .byteenable
		.cpu_data_master_read                                      (cpu_data_master_read),                                                //                                                    .read
		.cpu_data_master_readdata                                  (cpu_data_master_readdata),                                            //                                                    .readdata
		.cpu_data_master_write                                     (cpu_data_master_write),                                               //                                                    .write
		.cpu_data_master_writedata                                 (cpu_data_master_writedata),                                           //                                                    .writedata
		.cpu_data_master_debugaccess                               (cpu_data_master_debugaccess),                                         //                                                    .debugaccess
		.cpu_instruction_master_address                            (cpu_instruction_master_address),                                      //                              cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                        (cpu_instruction_master_waitrequest),                                  //                                                    .waitrequest
		.cpu_instruction_master_read                               (cpu_instruction_master_read),                                         //                                                    .read
		.cpu_instruction_master_readdata                           (cpu_instruction_master_readdata),                                     //                                                    .readdata
		.cpu_debug_mem_slave_address                               (mm_interconnect_0_cpu_debug_mem_slave_address),                       //                                 cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                 (mm_interconnect_0_cpu_debug_mem_slave_write),                         //                                                    .write
		.cpu_debug_mem_slave_read                                  (mm_interconnect_0_cpu_debug_mem_slave_read),                          //                                                    .read
		.cpu_debug_mem_slave_readdata                              (mm_interconnect_0_cpu_debug_mem_slave_readdata),                      //                                                    .readdata
		.cpu_debug_mem_slave_writedata                             (mm_interconnect_0_cpu_debug_mem_slave_writedata),                     //                                                    .writedata
		.cpu_debug_mem_slave_byteenable                            (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                    //                                                    .byteenable
		.cpu_debug_mem_slave_waitrequest                           (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                   //                                                    .waitrequest
		.cpu_debug_mem_slave_debugaccess                           (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                   //                                                    .debugaccess
		.div_freq_s1_address                                       (mm_interconnect_0_div_freq_s1_address),                               //                                         div_freq_s1.address
		.div_freq_s1_write                                         (mm_interconnect_0_div_freq_s1_write),                                 //                                                    .write
		.div_freq_s1_readdata                                      (mm_interconnect_0_div_freq_s1_readdata),                              //                                                    .readdata
		.div_freq_s1_writedata                                     (mm_interconnect_0_div_freq_s1_writedata),                             //                                                    .writedata
		.div_freq_s1_chipselect                                    (mm_interconnect_0_div_freq_s1_chipselect),                            //                                                    .chipselect
		.jtag_uart_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),               //                         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                 //                                                    .write
		.jtag_uart_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                  //                                                    .read
		.jtag_uart_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),              //                                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),             //                                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),           //                                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),            //                                                    .chipselect
		.leds_s1_address                                           (mm_interconnect_0_leds_s1_address),                                   //                                             leds_s1.address
		.leds_s1_write                                             (mm_interconnect_0_leds_s1_write),                                     //                                                    .write
		.leds_s1_readdata                                          (mm_interconnect_0_leds_s1_readdata),                                  //                                                    .readdata
		.leds_s1_writedata                                         (mm_interconnect_0_leds_s1_writedata),                                 //                                                    .writedata
		.leds_s1_chipselect                                        (mm_interconnect_0_leds_s1_chipselect),                                //                                                    .chipselect
		.noise_s1_address                                          (mm_interconnect_0_noise_s1_address),                                  //                                            noise_s1.address
		.noise_s1_write                                            (mm_interconnect_0_noise_s1_write),                                    //                                                    .write
		.noise_s1_readdata                                         (mm_interconnect_0_noise_s1_readdata),                                 //                                                    .readdata
		.noise_s1_writedata                                        (mm_interconnect_0_noise_s1_writedata),                                //                                                    .writedata
		.noise_s1_chipselect                                       (mm_interconnect_0_noise_s1_chipselect),                               //                                                    .chipselect
		.noise_en_s1_address                                       (mm_interconnect_0_noise_en_s1_address),                               //                                         noise_en_s1.address
		.noise_en_s1_write                                         (mm_interconnect_0_noise_en_s1_write),                                 //                                                    .write
		.noise_en_s1_readdata                                      (mm_interconnect_0_noise_en_s1_readdata),                              //                                                    .readdata
		.noise_en_s1_writedata                                     (mm_interconnect_0_noise_en_s1_writedata),                             //                                                    .writedata
		.noise_en_s1_chipselect                                    (mm_interconnect_0_noise_en_s1_chipselect),                            //                                                    .chipselect
		.noise_pulse_s1_address                                    (mm_interconnect_0_noise_pulse_s1_address),                            //                                      noise_pulse_s1.address
		.noise_pulse_s1_write                                      (mm_interconnect_0_noise_pulse_s1_write),                              //                                                    .write
		.noise_pulse_s1_readdata                                   (mm_interconnect_0_noise_pulse_s1_readdata),                           //                                                    .readdata
		.noise_pulse_s1_writedata                                  (mm_interconnect_0_noise_pulse_s1_writedata),                          //                                                    .writedata
		.noise_pulse_s1_chipselect                                 (mm_interconnect_0_noise_pulse_s1_chipselect),                         //                                                    .chipselect
		.RAM_jesus_s1_address                                      (mm_interconnect_0_ram_jesus_s1_address),                              //                                        RAM_jesus_s1.address
		.RAM_jesus_s1_write                                        (mm_interconnect_0_ram_jesus_s1_write),                                //                                                    .write
		.RAM_jesus_s1_readdata                                     (mm_interconnect_0_ram_jesus_s1_readdata),                             //                                                    .readdata
		.RAM_jesus_s1_writedata                                    (mm_interconnect_0_ram_jesus_s1_writedata),                            //                                                    .writedata
		.RAM_jesus_s1_byteenable                                   (mm_interconnect_0_ram_jesus_s1_byteenable),                           //                                                    .byteenable
		.RAM_jesus_s1_chipselect                                   (mm_interconnect_0_ram_jesus_s1_chipselect),                           //                                                    .chipselect
		.RAM_jesus_s1_clken                                        (mm_interconnect_0_ram_jesus_s1_clken),                                //                                                    .clken
		.sel_nota_s1_address                                       (mm_interconnect_0_sel_nota_s1_address),                               //                                         sel_nota_s1.address
		.sel_nota_s1_write                                         (mm_interconnect_0_sel_nota_s1_write),                                 //                                                    .write
		.sel_nota_s1_readdata                                      (mm_interconnect_0_sel_nota_s1_readdata),                              //                                                    .readdata
		.sel_nota_s1_writedata                                     (mm_interconnect_0_sel_nota_s1_writedata),                             //                                                    .writedata
		.sel_nota_s1_chipselect                                    (mm_interconnect_0_sel_nota_s1_chipselect),                            //                                                    .chipselect
		.sw_s1_address                                             (mm_interconnect_0_sw_s1_address),                                     //                                               sw_s1.address
		.sw_s1_readdata                                            (mm_interconnect_0_sw_s1_readdata),                                    //                                                    .readdata
		.sys_clk_s1_address                                        (mm_interconnect_0_sys_clk_s1_address),                                //                                          sys_clk_s1.address
		.sys_clk_s1_write                                          (mm_interconnect_0_sys_clk_s1_write),                                  //                                                    .write
		.sys_clk_s1_readdata                                       (mm_interconnect_0_sys_clk_s1_readdata),                               //                                                    .readdata
		.sys_clk_s1_writedata                                      (mm_interconnect_0_sys_clk_s1_writedata),                              //                                                    .writedata
		.sys_clk_s1_chipselect                                     (mm_interconnect_0_sys_clk_s1_chipselect),                             //                                                    .chipselect
		.timer_ece10243upb2016_0_avalon_slave_0_address            (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_address),    //              timer_ece10243upb2016_0_avalon_slave_0.address
		.timer_ece10243upb2016_0_avalon_slave_0_write              (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_write),      //                                                    .write
		.timer_ece10243upb2016_0_avalon_slave_0_readdata           (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_readdata),   //                                                    .readdata
		.timer_ece10243upb2016_0_avalon_slave_0_writedata          (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_writedata),  //                                                    .writedata
		.timer_ece10243upb2016_0_avalon_slave_0_chipselect         (mm_interconnect_0_timer_ece10243upb2016_0_avalon_slave_0_chipselect), //                                                    .chipselect
		.uart_s1_address                                           (mm_interconnect_0_uart_s1_address),                                   //                                             uart_s1.address
		.uart_s1_write                                             (mm_interconnect_0_uart_s1_write),                                     //                                                    .write
		.uart_s1_read                                              (mm_interconnect_0_uart_s1_read),                                      //                                                    .read
		.uart_s1_readdata                                          (mm_interconnect_0_uart_s1_readdata),                                  //                                                    .readdata
		.uart_s1_writedata                                         (mm_interconnect_0_uart_s1_writedata),                                 //                                                    .writedata
		.uart_s1_begintransfer                                     (mm_interconnect_0_uart_s1_begintransfer),                             //                                                    .begintransfer
		.uart_s1_chipselect                                        (mm_interconnect_0_uart_s1_chipselect)                                 //                                                    .chipselect
	);

	nios_practica_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
